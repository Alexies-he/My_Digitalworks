package fifo_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  `include "./fifo_sequence_item.sv"
endpackage 
