module fall_adder_down (
    input x,y,in,
    output out_in,out
);
    assign {out_in,out}=x+y+in;
endmodule