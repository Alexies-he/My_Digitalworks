`timescale 1ns/1ns
module tb_Ramdom_creater;
reg load,clk;
reg [4:0]D;//申明输入信号
wire out;//申明输出信号
initial 
	begin
	$display("start a clock pulse");
    $dumpfile("tb_Ramdom_creater.vcd");
    $dumpvars(0,tb_Ramdom_creater);
clk=0;load=0;D=5'b00001;//输入信号的波形
#10
clk=1;load=0;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
clk=0;load=1;D=5'b00001;
#10
clk=1;load=1;D=5'b00001;
#10
$stop;
$finish;
    end
    ramdom_creater U1(.clk(clk),.load(load),.D(D[2:0]),.out(out));
endmodule